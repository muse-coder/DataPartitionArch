VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO Ram_256_words
   CLASS BLOCK ;
   SIZE 229.045 BY 138.785 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  27.485 1.105 27.62 1.24 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  30.345 1.105 30.48 1.24 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.205 1.105 33.34 1.24 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.065 1.105 36.2 1.24 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.925 1.105 39.06 1.24 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.785 1.105 41.92 1.24 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.645 1.105 44.78 1.24 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.505 1.105 47.64 1.24 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.365 1.105 50.5 1.24 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.225 1.105 53.36 1.24 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.085 1.105 56.22 1.24 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.945 1.105 59.08 1.24 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.805 1.105 61.94 1.24 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.665 1.105 64.8 1.24 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.525 1.105 67.66 1.24 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.385 1.105 70.52 1.24 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.245 1.105 73.38 1.24 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.105 1.105 76.24 1.24 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.965 1.105 79.1 1.24 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.825 1.105 81.96 1.24 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.685 1.105 84.82 1.24 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.545 1.105 87.68 1.24 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.405 1.105 90.54 1.24 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.265 1.105 93.4 1.24 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.125 1.105 96.26 1.24 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.985 1.105 99.12 1.24 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.845 1.105 101.98 1.24 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.705 1.105 104.84 1.24 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.565 1.105 107.7 1.24 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.425 1.105 110.56 1.24 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.285 1.105 113.42 1.24 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.145 1.105 116.28 1.24 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  21.765 1.105 21.9 1.24 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24.625 1.105 24.76 1.24 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  16.045 48.6 16.18 48.735 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  16.045 51.33 16.18 51.465 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  16.045 53.54 16.18 53.675 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  16.045 56.27 16.18 56.405 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  16.045 58.48 16.18 58.615 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  16.045 61.21 16.18 61.345 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.145 137.545 204.28 137.68 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.285 137.545 201.42 137.68 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.725 22.47 212.86 22.605 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.725 19.74 212.86 19.875 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.725 17.53 212.86 17.665 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.725 14.8 212.86 14.935 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.725 12.59 212.86 12.725 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.725 9.86 212.86 9.995 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 4.01 0.42 4.145 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.625 136.17 228.76 136.305 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.2475 4.095 6.3825 4.23 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  222.5225 136.085 222.6575 136.22 ;
      END
   END clk1
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.1225 132.6775 39.2575 132.8125 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.8225 132.6775 43.9575 132.8125 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.5225 132.6775 48.6575 132.8125 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.2225 132.6775 53.3575 132.8125 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.9225 132.6775 58.0575 132.8125 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.6225 132.6775 62.7575 132.8125 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.3225 132.6775 67.4575 132.8125 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.0225 132.6775 72.1575 132.8125 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.7225 132.6775 76.8575 132.8125 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.4225 132.6775 81.5575 132.8125 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.1225 132.6775 86.2575 132.8125 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.8225 132.6775 90.9575 132.8125 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.5225 132.6775 95.6575 132.8125 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.2225 132.6775 100.3575 132.8125 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.9225 132.6775 105.0575 132.8125 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.6225 132.6775 109.7575 132.8125 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.3225 132.6775 114.4575 132.8125 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.0225 132.6775 119.1575 132.8125 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.7225 132.6775 123.8575 132.8125 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.4225 132.6775 128.5575 132.8125 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.1225 132.6775 133.2575 132.8125 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.8225 132.6775 137.9575 132.8125 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.5225 132.6775 142.6575 132.8125 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.2225 132.6775 147.3575 132.8125 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.9225 132.6775 152.0575 132.8125 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.6225 132.6775 156.7575 132.8125 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.3225 132.6775 161.4575 132.8125 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.0225 132.6775 166.1575 132.8125 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.7225 132.6775 170.8575 132.8125 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.4225 132.6775 175.5575 132.8125 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.1225 132.6775 180.2575 132.8125 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.8225 132.6775 184.9575 132.8125 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  21.8625 25.07 21.9975 25.205 ;
         LAYER metal3 ;
         RECT  35.9375 19.7075 189.6225 19.7775 ;
         LAYER metal3 ;
         RECT  35.9375 123.0075 190.7975 123.0775 ;
         LAYER metal3 ;
         RECT  21.8625 34.04 21.9975 34.175 ;
         LAYER metal3 ;
         RECT  200.54 119.9625 200.675 120.0975 ;
         LAYER metal3 ;
         RECT  34.7925 22.08 34.9275 22.215 ;
         LAYER metal3 ;
         RECT  95.8425 2.47 95.9775 2.605 ;
         LAYER metal4 ;
         RECT  193.78 23.5725 193.92 119.3925 ;
         LAYER metal4 ;
         RECT  228.2175 105.1625 228.3575 127.565 ;
         LAYER metal3 ;
         RECT  206.7125 37.03 206.8475 37.165 ;
         LAYER metal3 ;
         RECT  50.0825 2.47 50.2175 2.605 ;
         LAYER metal3 ;
         RECT  206.7125 34.04 206.8475 34.175 ;
         LAYER metal4 ;
         RECT  25.57 7.365 25.71 17.385 ;
         LAYER metal4 ;
         RECT  213.005 8.7525 213.145 23.7125 ;
         LAYER metal3 ;
         RECT  204.4275 136.18 204.5625 136.315 ;
         LAYER metal3 ;
         RECT  2.425 5.375 2.56 5.51 ;
         LAYER metal3 ;
         RECT  206.7125 43.01 206.8475 43.145 ;
         LAYER metal3 ;
         RECT  27.2025 2.47 27.3375 2.605 ;
         LAYER metal4 ;
         RECT  34.79 23.5725 34.93 119.3925 ;
         LAYER metal3 ;
         RECT  226.485 134.805 226.62 134.94 ;
         LAYER metal3 ;
         RECT  72.9625 2.47 73.0975 2.605 ;
         LAYER metal3 ;
         RECT  28.035 22.8675 28.17 23.0025 ;
         LAYER metal3 ;
         RECT  84.4025 2.47 84.5375 2.605 ;
         LAYER metal4 ;
         RECT  201.155 23.5725 201.295 119.4625 ;
         LAYER metal3 ;
         RECT  21.8625 37.03 21.9975 37.165 ;
         LAYER metal3 ;
         RECT  21.4825 2.47 21.6175 2.605 ;
         LAYER metal4 ;
         RECT  0.6875 12.75 0.8275 35.1525 ;
         LAYER metal3 ;
         RECT  61.5225 2.47 61.6575 2.605 ;
         LAYER metal3 ;
         RECT  193.7825 120.75 193.9175 120.885 ;
         LAYER metal3 ;
         RECT  35.9375 11.0575 185.6275 11.1275 ;
         LAYER metal3 ;
         RECT  21.8625 43.01 21.9975 43.145 ;
         LAYER metal3 ;
         RECT  206.7125 28.06 206.8475 28.195 ;
         LAYER metal4 ;
         RECT  27.415 23.5725 27.555 119.4625 ;
         LAYER metal3 ;
         RECT  21.8625 28.06 21.9975 28.195 ;
         LAYER metal4 ;
         RECT  203.0 125.4 203.14 135.42 ;
         LAYER metal3 ;
         RECT  21.8625 46.0 21.9975 46.135 ;
         LAYER metal4 ;
         RECT  18.48 5.3725 18.62 20.3325 ;
         LAYER metal3 ;
         RECT  206.7125 46.0 206.8475 46.135 ;
         LAYER metal4 ;
         RECT  192.7 20.4025 192.84 122.3125 ;
         LAYER metal4 ;
         RECT  210.285 124.9225 210.425 134.9425 ;
         LAYER metal3 ;
         RECT  206.7125 25.07 206.8475 25.205 ;
         LAYER metal4 ;
         RECT  15.76 47.4925 15.9 62.4525 ;
         LAYER metal3 ;
         RECT  107.2825 2.47 107.4175 2.605 ;
         LAYER metal3 ;
         RECT  38.6425 2.47 38.7775 2.605 ;
         LAYER metal3 ;
         RECT  35.9375 130.12 185.6275 130.19 ;
         LAYER metal4 ;
         RECT  35.87 20.4025 36.01 122.3125 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  192.24 20.4025 192.38 122.3125 ;
         LAYER metal3 ;
         RECT  20.335 35.535 20.47 35.67 ;
         LAYER metal4 ;
         RECT  25.48 23.54 25.62 119.4625 ;
         LAYER metal3 ;
         RECT  208.24 38.525 208.375 38.66 ;
         LAYER metal4 ;
         RECT  226.155 105.13 226.295 127.5325 ;
         LAYER metal3 ;
         RECT  110.1425 0.0 110.2775 0.135 ;
         LAYER metal3 ;
         RECT  208.24 47.495 208.375 47.63 ;
         LAYER metal3 ;
         RECT  208.24 32.545 208.375 32.68 ;
         LAYER metal3 ;
         RECT  35.9375 13.1075 185.6275 13.1775 ;
         LAYER metal4 ;
         RECT  18.62 47.4275 18.76 62.5175 ;
         LAYER metal3 ;
         RECT  30.0625 0.0 30.1975 0.135 ;
         LAYER metal3 ;
         RECT  87.2625 0.0 87.3975 0.135 ;
         LAYER metal3 ;
         RECT  41.5025 0.0 41.6375 0.135 ;
         LAYER metal3 ;
         RECT  208.24 35.535 208.375 35.67 ;
         LAYER metal3 ;
         RECT  20.335 47.495 20.47 47.63 ;
         LAYER metal4 ;
         RECT  204.6625 125.3325 204.8025 135.4875 ;
         LAYER metal3 ;
         RECT  98.7025 0.0 98.8375 0.135 ;
         LAYER metal3 ;
         RECT  208.24 26.565 208.375 26.7 ;
         LAYER metal3 ;
         RECT  24.3425 0.0 24.4775 0.135 ;
         LAYER metal4 ;
         RECT  210.145 8.6875 210.285 23.7775 ;
         LAYER metal3 ;
         RECT  35.9375 128.2275 185.6625 128.2975 ;
         LAYER metal3 ;
         RECT  20.335 32.545 20.47 32.68 ;
         LAYER metal3 ;
         RECT  208.24 23.575 208.375 23.71 ;
         LAYER metal3 ;
         RECT  20.335 38.525 20.47 38.66 ;
         LAYER metal3 ;
         RECT  208.24 29.555 208.375 29.69 ;
         LAYER metal3 ;
         RECT  75.8225 0.0 75.9575 0.135 ;
         LAYER metal3 ;
         RECT  20.335 29.555 20.47 29.69 ;
         LAYER metal3 ;
         RECT  201.5675 138.65 201.7025 138.785 ;
         LAYER metal3 ;
         RECT  208.24 41.515 208.375 41.65 ;
         LAYER metal4 ;
         RECT  200.595 23.54 200.735 119.425 ;
         LAYER metal3 ;
         RECT  35.9375 125.6275 189.655 125.6975 ;
         LAYER metal4 ;
         RECT  36.33 20.4025 36.47 122.3125 ;
         LAYER metal3 ;
         RECT  2.425 2.905 2.56 3.04 ;
         LAYER metal3 ;
         RECT  52.9425 0.0 53.0775 0.135 ;
         LAYER metal3 ;
         RECT  20.335 44.505 20.47 44.64 ;
         LAYER metal4 ;
         RECT  27.975 23.54 28.115 119.425 ;
         LAYER metal4 ;
         RECT  222.66 122.4525 222.8 137.4125 ;
         LAYER metal4 ;
         RECT  203.09 23.54 203.23 119.4625 ;
         LAYER metal4 ;
         RECT  23.9075 7.2975 24.0475 17.4525 ;
         LAYER metal4 ;
         RECT  6.105 2.9025 6.245 17.8625 ;
         LAYER metal3 ;
         RECT  20.335 41.515 20.47 41.65 ;
         LAYER metal3 ;
         RECT  208.24 44.505 208.375 44.64 ;
         LAYER metal3 ;
         RECT  35.9375 17.0875 189.655 17.1575 ;
         LAYER metal4 ;
         RECT  2.75 12.7825 2.89 35.185 ;
         LAYER metal3 ;
         RECT  226.485 137.275 226.62 137.41 ;
         LAYER metal3 ;
         RECT  20.335 23.575 20.47 23.71 ;
         LAYER metal3 ;
         RECT  20.335 26.565 20.47 26.7 ;
         LAYER metal3 ;
         RECT  64.3825 0.0 64.5175 0.135 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 228.905 138.645 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 228.905 138.645 ;
   LAYER  metal3 ;
      RECT  27.345 0.14 27.76 0.965 ;
      RECT  27.76 0.965 30.205 1.38 ;
      RECT  30.62 0.965 33.065 1.38 ;
      RECT  33.48 0.965 35.925 1.38 ;
      RECT  36.34 0.965 38.785 1.38 ;
      RECT  39.2 0.965 41.645 1.38 ;
      RECT  42.06 0.965 44.505 1.38 ;
      RECT  44.92 0.965 47.365 1.38 ;
      RECT  47.78 0.965 50.225 1.38 ;
      RECT  50.64 0.965 53.085 1.38 ;
      RECT  53.5 0.965 55.945 1.38 ;
      RECT  56.36 0.965 58.805 1.38 ;
      RECT  59.22 0.965 61.665 1.38 ;
      RECT  62.08 0.965 64.525 1.38 ;
      RECT  64.94 0.965 67.385 1.38 ;
      RECT  67.8 0.965 70.245 1.38 ;
      RECT  70.66 0.965 73.105 1.38 ;
      RECT  73.52 0.965 75.965 1.38 ;
      RECT  76.38 0.965 78.825 1.38 ;
      RECT  79.24 0.965 81.685 1.38 ;
      RECT  82.1 0.965 84.545 1.38 ;
      RECT  84.96 0.965 87.405 1.38 ;
      RECT  87.82 0.965 90.265 1.38 ;
      RECT  90.68 0.965 93.125 1.38 ;
      RECT  93.54 0.965 95.985 1.38 ;
      RECT  96.4 0.965 98.845 1.38 ;
      RECT  99.26 0.965 101.705 1.38 ;
      RECT  102.12 0.965 104.565 1.38 ;
      RECT  104.98 0.965 107.425 1.38 ;
      RECT  107.84 0.965 110.285 1.38 ;
      RECT  110.7 0.965 113.145 1.38 ;
      RECT  113.56 0.965 116.005 1.38 ;
      RECT  116.42 0.965 228.905 1.38 ;
      RECT  0.14 0.965 21.625 1.38 ;
      RECT  22.04 0.965 24.485 1.38 ;
      RECT  24.9 0.965 27.345 1.38 ;
      RECT  0.14 48.46 15.905 48.875 ;
      RECT  0.14 48.875 15.905 138.645 ;
      RECT  15.905 1.38 16.32 48.46 ;
      RECT  16.32 48.46 27.345 48.875 ;
      RECT  16.32 48.875 27.345 138.645 ;
      RECT  15.905 48.875 16.32 51.19 ;
      RECT  15.905 51.605 16.32 53.4 ;
      RECT  15.905 53.815 16.32 56.13 ;
      RECT  15.905 56.545 16.32 58.34 ;
      RECT  15.905 58.755 16.32 61.07 ;
      RECT  15.905 61.485 16.32 138.645 ;
      RECT  204.005 137.82 204.42 138.645 ;
      RECT  204.42 137.82 228.905 138.645 ;
      RECT  27.76 137.405 201.145 137.82 ;
      RECT  201.56 137.405 204.005 137.82 ;
      RECT  204.42 1.38 212.585 22.33 ;
      RECT  204.42 22.33 212.585 22.745 ;
      RECT  212.585 22.745 213.0 137.405 ;
      RECT  213.0 1.38 228.905 22.33 ;
      RECT  213.0 22.33 228.905 22.745 ;
      RECT  212.585 20.015 213.0 22.33 ;
      RECT  212.585 17.805 213.0 19.6 ;
      RECT  212.585 15.075 213.0 17.39 ;
      RECT  212.585 12.865 213.0 14.66 ;
      RECT  212.585 1.38 213.0 9.72 ;
      RECT  212.585 10.135 213.0 12.45 ;
      RECT  0.14 1.38 0.145 3.87 ;
      RECT  0.14 3.87 0.145 4.285 ;
      RECT  0.14 4.285 0.145 48.46 ;
      RECT  0.145 1.38 0.56 3.87 ;
      RECT  0.145 4.285 0.56 48.46 ;
      RECT  228.485 22.745 228.9 136.03 ;
      RECT  228.485 136.445 228.9 137.405 ;
      RECT  228.9 22.745 228.905 136.03 ;
      RECT  228.9 136.03 228.905 136.445 ;
      RECT  228.9 136.445 228.905 137.405 ;
      RECT  0.56 3.87 6.1075 3.955 ;
      RECT  0.56 3.955 6.1075 4.285 ;
      RECT  6.1075 3.87 6.5225 3.955 ;
      RECT  6.5225 3.87 15.905 3.955 ;
      RECT  6.5225 3.955 15.905 4.285 ;
      RECT  0.56 4.285 6.1075 4.37 ;
      RECT  6.1075 4.37 6.5225 48.46 ;
      RECT  6.5225 4.285 15.905 4.37 ;
      RECT  6.5225 4.37 15.905 48.46 ;
      RECT  213.0 22.745 222.3825 135.945 ;
      RECT  213.0 135.945 222.3825 136.03 ;
      RECT  222.3825 22.745 222.7975 135.945 ;
      RECT  222.7975 135.945 228.485 136.03 ;
      RECT  213.0 136.03 222.3825 136.36 ;
      RECT  213.0 136.36 222.3825 136.445 ;
      RECT  222.3825 136.36 222.7975 136.445 ;
      RECT  222.7975 136.03 228.485 136.36 ;
      RECT  222.7975 136.36 228.485 136.445 ;
      RECT  27.76 132.5375 38.9825 132.9525 ;
      RECT  27.76 132.9525 38.9825 137.405 ;
      RECT  38.9825 132.9525 39.3975 137.405 ;
      RECT  39.3975 132.9525 204.005 137.405 ;
      RECT  39.3975 132.5375 43.6825 132.9525 ;
      RECT  44.0975 132.5375 48.3825 132.9525 ;
      RECT  48.7975 132.5375 53.0825 132.9525 ;
      RECT  53.4975 132.5375 57.7825 132.9525 ;
      RECT  58.1975 132.5375 62.4825 132.9525 ;
      RECT  62.8975 132.5375 67.1825 132.9525 ;
      RECT  67.5975 132.5375 71.8825 132.9525 ;
      RECT  72.2975 132.5375 76.5825 132.9525 ;
      RECT  76.9975 132.5375 81.2825 132.9525 ;
      RECT  81.6975 132.5375 85.9825 132.9525 ;
      RECT  86.3975 132.5375 90.6825 132.9525 ;
      RECT  91.0975 132.5375 95.3825 132.9525 ;
      RECT  95.7975 132.5375 100.0825 132.9525 ;
      RECT  100.4975 132.5375 104.7825 132.9525 ;
      RECT  105.1975 132.5375 109.4825 132.9525 ;
      RECT  109.8975 132.5375 114.1825 132.9525 ;
      RECT  114.5975 132.5375 118.8825 132.9525 ;
      RECT  119.2975 132.5375 123.5825 132.9525 ;
      RECT  123.9975 132.5375 128.2825 132.9525 ;
      RECT  128.6975 132.5375 132.9825 132.9525 ;
      RECT  133.3975 132.5375 137.6825 132.9525 ;
      RECT  138.0975 132.5375 142.3825 132.9525 ;
      RECT  142.7975 132.5375 147.0825 132.9525 ;
      RECT  147.4975 132.5375 151.7825 132.9525 ;
      RECT  152.1975 132.5375 156.4825 132.9525 ;
      RECT  156.8975 132.5375 161.1825 132.9525 ;
      RECT  161.5975 132.5375 165.8825 132.9525 ;
      RECT  166.2975 132.5375 170.5825 132.9525 ;
      RECT  170.9975 132.5375 175.2825 132.9525 ;
      RECT  175.6975 132.5375 179.9825 132.9525 ;
      RECT  180.3975 132.5375 184.6825 132.9525 ;
      RECT  185.0975 132.5375 204.005 132.9525 ;
      RECT  16.32 24.93 21.7225 25.345 ;
      RECT  22.1375 24.93 27.345 25.345 ;
      RECT  22.1375 25.345 27.345 48.46 ;
      RECT  27.76 1.38 35.7975 19.5675 ;
      RECT  27.76 19.5675 35.7975 19.9175 ;
      RECT  189.7625 19.5675 204.005 19.9175 ;
      RECT  35.7975 19.9175 38.9825 122.8675 ;
      RECT  38.9825 19.9175 39.3975 122.8675 ;
      RECT  39.3975 19.9175 189.7625 122.8675 ;
      RECT  189.7625 19.9175 190.9375 122.8675 ;
      RECT  190.9375 122.8675 204.005 123.2175 ;
      RECT  190.9375 123.2175 204.005 132.5375 ;
      RECT  190.9375 19.9175 200.4 119.8225 ;
      RECT  190.9375 119.8225 200.4 120.2375 ;
      RECT  200.4 19.9175 200.815 119.8225 ;
      RECT  200.4 120.2375 200.815 122.8675 ;
      RECT  200.815 19.9175 204.005 119.8225 ;
      RECT  200.815 119.8225 204.005 120.2375 ;
      RECT  200.815 120.2375 204.005 122.8675 ;
      RECT  27.76 19.9175 34.6525 21.94 ;
      RECT  27.76 21.94 34.6525 22.355 ;
      RECT  34.6525 19.9175 35.0675 21.94 ;
      RECT  34.6525 22.355 35.0675 132.5375 ;
      RECT  35.0675 19.9175 35.7975 21.94 ;
      RECT  35.0675 21.94 35.7975 22.355 ;
      RECT  35.0675 22.355 35.7975 132.5375 ;
      RECT  39.3975 1.38 95.7025 2.33 ;
      RECT  95.7025 1.38 96.1175 2.33 ;
      RECT  96.1175 1.38 189.7625 2.33 ;
      RECT  204.42 22.745 206.5725 36.89 ;
      RECT  204.42 36.89 206.5725 37.305 ;
      RECT  206.9875 36.89 212.585 37.305 ;
      RECT  39.3975 2.33 49.9425 2.745 ;
      RECT  206.5725 34.315 206.9875 36.89 ;
      RECT  204.005 1.38 204.2875 136.04 ;
      RECT  204.005 136.04 204.2875 136.455 ;
      RECT  204.005 136.455 204.2875 137.405 ;
      RECT  204.2875 1.38 204.42 136.04 ;
      RECT  204.2875 136.455 204.42 137.405 ;
      RECT  204.42 37.305 204.7025 136.04 ;
      RECT  204.42 136.455 204.7025 137.405 ;
      RECT  204.7025 37.305 206.5725 136.04 ;
      RECT  204.7025 136.04 206.5725 136.455 ;
      RECT  204.7025 136.455 206.5725 137.405 ;
      RECT  0.56 4.37 2.285 5.235 ;
      RECT  0.56 5.235 2.285 5.65 ;
      RECT  0.56 5.65 2.285 48.46 ;
      RECT  2.285 4.37 2.7 5.235 ;
      RECT  2.285 5.65 2.7 48.46 ;
      RECT  2.7 4.37 6.1075 5.235 ;
      RECT  2.7 5.235 6.1075 5.65 ;
      RECT  2.7 5.65 6.1075 48.46 ;
      RECT  206.5725 37.305 206.9875 42.87 ;
      RECT  27.345 1.38 27.4775 2.33 ;
      RECT  27.345 2.745 27.4775 138.645 ;
      RECT  27.4775 1.38 27.76 2.33 ;
      RECT  27.4775 2.33 27.76 2.745 ;
      RECT  27.4775 2.745 27.76 138.645 ;
      RECT  22.1375 1.38 27.0625 2.33 ;
      RECT  22.1375 2.33 27.0625 2.745 ;
      RECT  22.1375 2.745 27.0625 24.93 ;
      RECT  27.0625 1.38 27.345 2.33 ;
      RECT  27.0625 2.745 27.345 24.93 ;
      RECT  222.7975 22.745 226.345 134.665 ;
      RECT  222.7975 134.665 226.345 135.08 ;
      RECT  222.7975 135.08 226.345 135.945 ;
      RECT  226.345 22.745 226.76 134.665 ;
      RECT  226.345 135.08 226.76 135.945 ;
      RECT  226.76 22.745 228.485 134.665 ;
      RECT  226.76 134.665 228.485 135.08 ;
      RECT  226.76 135.08 228.485 135.945 ;
      RECT  27.76 22.355 27.895 22.7275 ;
      RECT  27.76 22.7275 27.895 23.1425 ;
      RECT  27.76 23.1425 27.895 132.5375 ;
      RECT  27.895 22.355 28.31 22.7275 ;
      RECT  27.895 23.1425 28.31 132.5375 ;
      RECT  28.31 22.355 34.6525 22.7275 ;
      RECT  28.31 22.7275 34.6525 23.1425 ;
      RECT  28.31 23.1425 34.6525 132.5375 ;
      RECT  73.2375 2.33 84.2625 2.745 ;
      RECT  84.6775 2.33 95.7025 2.745 ;
      RECT  21.7225 34.315 22.1375 36.89 ;
      RECT  16.32 1.38 21.3425 2.33 ;
      RECT  16.32 2.33 21.3425 2.745 ;
      RECT  21.3425 1.38 21.7225 2.33 ;
      RECT  21.3425 2.745 21.7225 24.93 ;
      RECT  21.7225 1.38 21.7575 2.33 ;
      RECT  21.7225 2.745 21.7575 24.93 ;
      RECT  21.7575 1.38 22.1375 2.33 ;
      RECT  21.7575 2.33 22.1375 2.745 ;
      RECT  21.7575 2.745 22.1375 24.93 ;
      RECT  50.3575 2.33 61.3825 2.745 ;
      RECT  61.7975 2.33 72.8225 2.745 ;
      RECT  190.9375 120.2375 193.6425 120.61 ;
      RECT  190.9375 120.61 193.6425 121.025 ;
      RECT  190.9375 121.025 193.6425 122.8675 ;
      RECT  193.6425 120.2375 194.0575 120.61 ;
      RECT  193.6425 121.025 194.0575 122.8675 ;
      RECT  194.0575 120.2375 200.4 120.61 ;
      RECT  194.0575 120.61 200.4 121.025 ;
      RECT  194.0575 121.025 200.4 122.8675 ;
      RECT  38.9825 1.38 39.3975 10.9175 ;
      RECT  39.3975 2.745 95.7025 10.9175 ;
      RECT  95.7025 2.745 96.1175 10.9175 ;
      RECT  96.1175 2.745 185.7675 10.9175 ;
      RECT  185.7675 2.745 189.7625 10.9175 ;
      RECT  185.7675 10.9175 189.7625 11.2675 ;
      RECT  21.7225 37.305 22.1375 42.87 ;
      RECT  206.5725 28.335 206.9875 33.9 ;
      RECT  21.7225 25.345 22.1375 27.92 ;
      RECT  21.7225 28.335 22.1375 33.9 ;
      RECT  21.7225 43.285 22.1375 45.86 ;
      RECT  21.7225 46.275 22.1375 48.46 ;
      RECT  206.5725 43.285 206.9875 45.86 ;
      RECT  206.5725 46.275 206.9875 137.405 ;
      RECT  206.5725 22.745 206.9875 24.93 ;
      RECT  206.5725 25.345 206.9875 27.92 ;
      RECT  96.1175 2.33 107.1425 2.745 ;
      RECT  107.5575 2.33 189.7625 2.745 ;
      RECT  35.7975 1.38 38.5025 2.33 ;
      RECT  35.7975 2.33 38.5025 2.745 ;
      RECT  35.7975 2.745 38.5025 10.9175 ;
      RECT  38.5025 1.38 38.9175 2.33 ;
      RECT  38.5025 2.745 38.9175 10.9175 ;
      RECT  38.9175 1.38 38.9825 2.33 ;
      RECT  38.9175 2.33 38.9825 2.745 ;
      RECT  38.9175 2.745 38.9825 10.9175 ;
      RECT  35.7975 130.33 38.9825 132.5375 ;
      RECT  38.9825 130.33 39.3975 132.5375 ;
      RECT  39.3975 130.33 185.7675 132.5375 ;
      RECT  185.7675 129.98 189.7625 130.33 ;
      RECT  185.7675 130.33 189.7625 132.5375 ;
      RECT  16.32 25.345 20.195 35.395 ;
      RECT  16.32 35.395 20.195 35.81 ;
      RECT  16.32 35.81 20.195 48.46 ;
      RECT  20.61 25.345 21.7225 35.395 ;
      RECT  20.61 35.395 21.7225 35.81 ;
      RECT  20.61 35.81 21.7225 48.46 ;
      RECT  206.9875 37.305 208.1 38.385 ;
      RECT  206.9875 38.385 208.1 38.8 ;
      RECT  206.9875 38.8 208.1 137.405 ;
      RECT  208.1 37.305 208.515 38.385 ;
      RECT  208.515 37.305 212.585 38.385 ;
      RECT  208.515 38.385 212.585 38.8 ;
      RECT  208.515 38.8 212.585 137.405 ;
      RECT  27.76 0.275 110.0025 0.965 ;
      RECT  110.0025 0.275 110.4175 0.965 ;
      RECT  110.4175 0.14 228.905 0.275 ;
      RECT  110.4175 0.275 228.905 0.965 ;
      RECT  208.1 47.77 208.515 137.405 ;
      RECT  206.9875 22.745 208.1 32.405 ;
      RECT  206.9875 32.405 208.1 32.82 ;
      RECT  206.9875 32.82 208.1 36.89 ;
      RECT  208.515 22.745 212.585 32.405 ;
      RECT  208.515 32.405 212.585 32.82 ;
      RECT  208.515 32.82 212.585 36.89 ;
      RECT  35.7975 11.2675 38.9825 12.9675 ;
      RECT  38.9825 11.2675 39.3975 12.9675 ;
      RECT  39.3975 11.2675 95.7025 12.9675 ;
      RECT  95.7025 11.2675 96.1175 12.9675 ;
      RECT  96.1175 11.2675 185.7675 12.9675 ;
      RECT  27.76 0.14 29.9225 0.275 ;
      RECT  30.3375 0.14 41.3625 0.275 ;
      RECT  208.1 32.82 208.515 35.395 ;
      RECT  208.1 35.81 208.515 36.89 ;
      RECT  20.195 47.77 20.61 48.46 ;
      RECT  87.5375 0.14 98.5625 0.275 ;
      RECT  98.9775 0.14 110.0025 0.275 ;
      RECT  0.14 0.14 24.2025 0.275 ;
      RECT  0.14 0.275 24.2025 0.965 ;
      RECT  24.2025 0.275 24.6175 0.965 ;
      RECT  24.6175 0.14 27.345 0.275 ;
      RECT  24.6175 0.275 27.345 0.965 ;
      RECT  35.7975 128.4375 38.9825 129.98 ;
      RECT  38.9825 128.4375 39.3975 129.98 ;
      RECT  39.3975 128.4375 185.7675 129.98 ;
      RECT  185.7675 128.4375 185.8025 129.98 ;
      RECT  185.8025 128.0875 189.7625 128.4375 ;
      RECT  185.8025 128.4375 189.7625 129.98 ;
      RECT  20.195 32.82 20.61 35.395 ;
      RECT  208.1 22.745 208.515 23.435 ;
      RECT  208.1 23.85 208.515 26.425 ;
      RECT  20.195 35.81 20.61 38.385 ;
      RECT  208.1 26.84 208.515 29.415 ;
      RECT  208.1 29.83 208.515 32.405 ;
      RECT  76.0975 0.14 87.1225 0.275 ;
      RECT  20.195 29.83 20.61 32.405 ;
      RECT  27.76 137.82 201.4275 138.51 ;
      RECT  27.76 138.51 201.4275 138.645 ;
      RECT  201.4275 137.82 201.8425 138.51 ;
      RECT  201.8425 137.82 204.005 138.51 ;
      RECT  201.8425 138.51 204.005 138.645 ;
      RECT  208.1 38.8 208.515 41.375 ;
      RECT  189.7625 123.2175 189.795 125.4875 ;
      RECT  189.7625 125.8375 189.795 132.5375 ;
      RECT  189.795 123.2175 190.9375 125.4875 ;
      RECT  189.795 125.4875 190.9375 125.8375 ;
      RECT  189.795 125.8375 190.9375 132.5375 ;
      RECT  35.7975 123.2175 38.9825 125.4875 ;
      RECT  35.7975 125.8375 38.9825 128.0875 ;
      RECT  38.9825 123.2175 39.3975 125.4875 ;
      RECT  38.9825 125.8375 39.3975 128.0875 ;
      RECT  39.3975 123.2175 185.7675 125.4875 ;
      RECT  39.3975 125.8375 185.7675 128.0875 ;
      RECT  185.7675 123.2175 185.8025 125.4875 ;
      RECT  185.7675 125.8375 185.8025 128.0875 ;
      RECT  185.8025 123.2175 189.7625 125.4875 ;
      RECT  185.8025 125.8375 189.7625 128.0875 ;
      RECT  0.56 1.38 2.285 2.765 ;
      RECT  0.56 2.765 2.285 3.18 ;
      RECT  0.56 3.18 2.285 3.87 ;
      RECT  2.285 1.38 2.7 2.765 ;
      RECT  2.285 3.18 2.7 3.87 ;
      RECT  2.7 1.38 15.905 2.765 ;
      RECT  2.7 2.765 15.905 3.18 ;
      RECT  2.7 3.18 15.905 3.87 ;
      RECT  41.7775 0.14 52.8025 0.275 ;
      RECT  20.195 44.78 20.61 47.355 ;
      RECT  20.195 38.8 20.61 41.375 ;
      RECT  20.195 41.79 20.61 44.365 ;
      RECT  208.1 41.79 208.515 44.365 ;
      RECT  208.1 44.78 208.515 47.355 ;
      RECT  189.7625 1.38 189.795 16.9475 ;
      RECT  189.7625 17.2975 189.795 19.5675 ;
      RECT  189.795 1.38 204.005 16.9475 ;
      RECT  189.795 16.9475 204.005 17.2975 ;
      RECT  189.795 17.2975 204.005 19.5675 ;
      RECT  185.7675 11.2675 189.7625 16.9475 ;
      RECT  185.7675 17.2975 189.7625 19.5675 ;
      RECT  35.7975 13.3175 38.9825 16.9475 ;
      RECT  35.7975 17.2975 38.9825 19.5675 ;
      RECT  38.9825 13.3175 39.3975 16.9475 ;
      RECT  38.9825 17.2975 39.3975 19.5675 ;
      RECT  39.3975 13.3175 95.7025 16.9475 ;
      RECT  39.3975 17.2975 95.7025 19.5675 ;
      RECT  95.7025 13.3175 96.1175 16.9475 ;
      RECT  95.7025 17.2975 96.1175 19.5675 ;
      RECT  96.1175 13.3175 185.7675 16.9475 ;
      RECT  96.1175 17.2975 185.7675 19.5675 ;
      RECT  204.42 137.405 226.345 137.55 ;
      RECT  204.42 137.55 226.345 137.82 ;
      RECT  226.345 137.55 226.76 137.82 ;
      RECT  226.76 137.405 228.905 137.55 ;
      RECT  226.76 137.55 228.905 137.82 ;
      RECT  213.0 136.445 226.345 137.135 ;
      RECT  213.0 137.135 226.345 137.405 ;
      RECT  226.345 136.445 226.76 137.135 ;
      RECT  226.76 136.445 228.485 137.135 ;
      RECT  226.76 137.135 228.485 137.405 ;
      RECT  16.32 2.745 20.195 23.435 ;
      RECT  16.32 23.435 20.195 23.85 ;
      RECT  16.32 23.85 20.195 24.93 ;
      RECT  20.195 2.745 20.61 23.435 ;
      RECT  20.195 23.85 20.61 24.93 ;
      RECT  20.61 2.745 21.3425 23.435 ;
      RECT  20.61 23.435 21.3425 23.85 ;
      RECT  20.61 23.85 21.3425 24.93 ;
      RECT  20.195 25.345 20.61 26.425 ;
      RECT  20.195 26.84 20.61 29.415 ;
      RECT  53.2175 0.14 64.2425 0.275 ;
      RECT  64.6575 0.14 75.6825 0.275 ;
   LAYER  metal4 ;
      RECT  193.5 0.14 194.2 23.2925 ;
      RECT  193.5 119.6725 194.2 138.645 ;
      RECT  227.9375 23.2925 228.6375 104.8825 ;
      RECT  228.6375 23.2925 228.905 104.8825 ;
      RECT  228.6375 104.8825 228.905 119.6725 ;
      RECT  227.9375 127.845 228.6375 138.645 ;
      RECT  228.6375 119.6725 228.905 127.845 ;
      RECT  228.6375 127.845 228.905 138.645 ;
      RECT  25.29 0.14 25.99 7.085 ;
      RECT  25.99 0.14 193.5 7.085 ;
      RECT  25.99 7.085 193.5 17.665 ;
      RECT  212.725 0.14 213.425 8.4725 ;
      RECT  213.425 0.14 228.905 8.4725 ;
      RECT  213.425 8.4725 228.905 23.2925 ;
      RECT  212.725 23.9925 213.425 104.8825 ;
      RECT  213.425 23.2925 227.9375 23.9925 ;
      RECT  194.2 119.7425 200.875 127.845 ;
      RECT  200.875 119.7425 201.575 127.845 ;
      RECT  0.14 7.085 0.4075 12.47 ;
      RECT  0.14 12.47 0.4075 17.665 ;
      RECT  0.4075 7.085 1.1075 12.47 ;
      RECT  0.14 17.665 0.4075 23.2925 ;
      RECT  0.14 23.2925 0.4075 35.4325 ;
      RECT  0.14 35.4325 0.4075 119.6725 ;
      RECT  0.4075 35.4325 1.1075 119.6725 ;
      RECT  0.14 119.7425 27.135 138.645 ;
      RECT  27.135 119.7425 27.835 138.645 ;
      RECT  194.2 127.845 202.72 135.7 ;
      RECT  194.2 135.7 202.72 138.645 ;
      RECT  202.72 135.7 203.42 138.645 ;
      RECT  201.575 119.7425 202.72 125.12 ;
      RECT  201.575 125.12 202.72 127.845 ;
      RECT  202.72 119.7425 203.42 125.12 ;
      RECT  18.2 0.14 18.9 5.0925 ;
      RECT  18.9 0.14 25.29 5.0925 ;
      RECT  18.2 20.6125 18.9 23.2925 ;
      RECT  25.99 17.665 192.42 20.1225 ;
      RECT  192.42 17.665 193.12 20.1225 ;
      RECT  193.12 17.665 193.5 20.1225 ;
      RECT  193.12 20.1225 193.5 23.2925 ;
      RECT  193.12 23.2925 193.5 119.6725 ;
      RECT  193.12 119.6725 193.5 119.7425 ;
      RECT  27.835 122.5925 192.42 138.645 ;
      RECT  192.42 122.5925 193.12 138.645 ;
      RECT  193.12 119.7425 193.5 122.5925 ;
      RECT  193.12 122.5925 193.5 138.645 ;
      RECT  210.005 135.2225 210.705 135.7 ;
      RECT  203.42 119.7425 210.005 124.6425 ;
      RECT  210.005 119.7425 210.705 124.6425 ;
      RECT  1.1075 47.2125 15.48 62.7325 ;
      RECT  1.1075 62.7325 15.48 119.6725 ;
      RECT  15.48 35.4325 16.18 47.2125 ;
      RECT  15.48 62.7325 16.18 119.6725 ;
      RECT  35.21 23.2925 35.59 119.6725 ;
      RECT  27.835 119.7425 35.59 122.5925 ;
      RECT  25.29 17.665 25.9 23.26 ;
      RECT  25.9 17.665 25.99 23.26 ;
      RECT  25.9 23.26 25.99 23.2925 ;
      RECT  0.14 119.6725 25.2 119.7425 ;
      RECT  25.9 119.6725 27.135 119.7425 ;
      RECT  25.9 23.2925 27.135 35.4325 ;
      RECT  18.9 20.6125 25.2 23.26 ;
      RECT  18.9 23.26 25.2 23.2925 ;
      RECT  25.2 20.6125 25.29 23.26 ;
      RECT  25.9 35.4325 27.135 47.2125 ;
      RECT  25.9 47.2125 27.135 62.7325 ;
      RECT  25.9 62.7325 27.135 119.6725 ;
      RECT  213.425 23.9925 225.875 104.85 ;
      RECT  213.425 104.85 225.875 104.8825 ;
      RECT  225.875 23.9925 226.575 104.85 ;
      RECT  226.575 23.9925 227.9375 104.85 ;
      RECT  226.575 104.85 227.9375 104.8825 ;
      RECT  226.575 104.8825 227.9375 119.6725 ;
      RECT  226.575 119.6725 227.9375 119.7425 ;
      RECT  226.575 119.7425 227.9375 124.6425 ;
      RECT  226.575 124.6425 227.9375 125.12 ;
      RECT  225.875 127.8125 226.575 127.845 ;
      RECT  226.575 125.12 227.9375 127.8125 ;
      RECT  226.575 127.8125 227.9375 127.845 ;
      RECT  16.18 35.4325 18.34 47.1475 ;
      RECT  16.18 47.1475 18.34 47.2125 ;
      RECT  18.34 35.4325 19.04 47.1475 ;
      RECT  19.04 35.4325 25.2 47.1475 ;
      RECT  19.04 47.1475 25.2 47.2125 ;
      RECT  16.18 47.2125 18.34 62.7325 ;
      RECT  19.04 47.2125 25.2 62.7325 ;
      RECT  16.18 62.7325 18.34 62.7975 ;
      RECT  16.18 62.7975 18.34 119.6725 ;
      RECT  18.34 62.7975 19.04 119.6725 ;
      RECT  19.04 62.7325 25.2 62.7975 ;
      RECT  19.04 62.7975 25.2 119.6725 ;
      RECT  203.42 135.7 204.3825 135.7675 ;
      RECT  203.42 135.7675 204.3825 138.645 ;
      RECT  204.3825 135.7675 205.0825 138.645 ;
      RECT  203.42 127.845 204.3825 135.2225 ;
      RECT  205.0825 127.845 210.005 135.2225 ;
      RECT  203.42 135.2225 204.3825 135.7 ;
      RECT  205.0825 135.2225 210.005 135.7 ;
      RECT  203.42 124.6425 204.3825 125.0525 ;
      RECT  203.42 125.0525 204.3825 125.12 ;
      RECT  204.3825 124.6425 205.0825 125.0525 ;
      RECT  205.0825 124.6425 210.005 125.0525 ;
      RECT  205.0825 125.0525 210.005 125.12 ;
      RECT  203.42 125.12 204.3825 127.845 ;
      RECT  205.0825 125.12 210.005 127.845 ;
      RECT  194.2 0.14 209.865 8.4075 ;
      RECT  194.2 8.4075 209.865 8.4725 ;
      RECT  209.865 0.14 210.565 8.4075 ;
      RECT  210.565 0.14 212.725 8.4075 ;
      RECT  210.565 8.4075 212.725 8.4725 ;
      RECT  210.565 8.4725 212.725 23.2925 ;
      RECT  210.565 23.2925 212.725 23.9925 ;
      RECT  209.865 24.0575 210.565 104.8825 ;
      RECT  210.565 23.9925 212.725 24.0575 ;
      RECT  210.565 24.0575 212.725 104.8825 ;
      RECT  194.2 104.8825 200.315 119.6725 ;
      RECT  194.2 119.6725 200.315 119.705 ;
      RECT  194.2 119.705 200.315 119.7425 ;
      RECT  200.315 119.705 200.875 119.7425 ;
      RECT  194.2 23.2925 200.315 23.9925 ;
      RECT  194.2 23.9925 200.315 104.8825 ;
      RECT  194.2 8.4725 200.315 23.26 ;
      RECT  194.2 23.26 200.315 23.2925 ;
      RECT  200.315 8.4725 201.015 23.26 ;
      RECT  201.015 8.4725 209.865 23.26 ;
      RECT  36.75 20.1225 191.96 23.2925 ;
      RECT  36.75 23.2925 191.96 119.6725 ;
      RECT  36.75 119.6725 191.96 119.7425 ;
      RECT  36.75 119.7425 191.96 122.5925 ;
      RECT  28.395 23.2925 34.51 35.4325 ;
      RECT  28.395 35.4325 34.51 119.6725 ;
      RECT  25.99 20.1225 27.695 23.26 ;
      RECT  25.99 23.26 27.695 23.2925 ;
      RECT  27.695 20.1225 28.395 23.26 ;
      RECT  28.395 20.1225 35.59 23.26 ;
      RECT  28.395 23.26 35.59 23.2925 ;
      RECT  27.835 119.705 28.395 119.7425 ;
      RECT  28.395 119.6725 35.59 119.705 ;
      RECT  28.395 119.705 35.59 119.7425 ;
      RECT  210.705 127.845 222.38 135.2225 ;
      RECT  223.08 127.845 227.9375 135.2225 ;
      RECT  210.705 135.2225 222.38 135.7 ;
      RECT  223.08 135.2225 227.9375 135.7 ;
      RECT  210.705 119.7425 222.38 122.1725 ;
      RECT  210.705 122.1725 222.38 124.6425 ;
      RECT  222.38 119.7425 223.08 122.1725 ;
      RECT  223.08 119.7425 225.875 122.1725 ;
      RECT  223.08 122.1725 225.875 124.6425 ;
      RECT  210.705 124.6425 222.38 125.12 ;
      RECT  223.08 124.6425 225.875 125.12 ;
      RECT  210.705 125.12 222.38 127.8125 ;
      RECT  223.08 125.12 225.875 127.8125 ;
      RECT  210.705 127.8125 222.38 127.845 ;
      RECT  223.08 127.8125 225.875 127.845 ;
      RECT  205.0825 135.7 222.38 135.7675 ;
      RECT  223.08 135.7 227.9375 135.7675 ;
      RECT  205.0825 135.7675 222.38 137.6925 ;
      RECT  205.0825 137.6925 222.38 138.645 ;
      RECT  222.38 137.6925 223.08 138.645 ;
      RECT  223.08 135.7675 227.9375 137.6925 ;
      RECT  223.08 137.6925 227.9375 138.645 ;
      RECT  201.575 104.8825 202.81 119.6725 ;
      RECT  203.51 104.8825 225.875 119.6725 ;
      RECT  201.575 119.6725 202.81 119.7425 ;
      RECT  203.51 119.6725 225.875 119.7425 ;
      RECT  201.575 23.2925 202.81 23.9925 ;
      RECT  203.51 23.2925 209.865 23.9925 ;
      RECT  201.575 23.9925 202.81 24.0575 ;
      RECT  203.51 23.9925 209.865 24.0575 ;
      RECT  201.575 24.0575 202.81 104.8825 ;
      RECT  203.51 24.0575 209.865 104.8825 ;
      RECT  201.015 23.26 202.81 23.2925 ;
      RECT  203.51 23.26 209.865 23.2925 ;
      RECT  18.9 5.0925 23.6275 7.0175 ;
      RECT  18.9 7.0175 23.6275 7.085 ;
      RECT  23.6275 5.0925 24.3275 7.0175 ;
      RECT  24.3275 5.0925 25.29 7.0175 ;
      RECT  24.3275 7.0175 25.29 7.085 ;
      RECT  18.9 7.085 23.6275 12.47 ;
      RECT  24.3275 7.085 25.29 12.47 ;
      RECT  18.9 12.47 23.6275 17.665 ;
      RECT  24.3275 12.47 25.29 17.665 ;
      RECT  18.9 17.665 23.6275 17.7325 ;
      RECT  18.9 17.7325 23.6275 20.6125 ;
      RECT  23.6275 17.7325 24.3275 20.6125 ;
      RECT  24.3275 17.665 25.29 17.7325 ;
      RECT  24.3275 17.7325 25.29 20.6125 ;
      RECT  0.14 0.14 5.825 2.6225 ;
      RECT  0.14 2.6225 5.825 5.0925 ;
      RECT  5.825 0.14 6.525 2.6225 ;
      RECT  6.525 0.14 18.2 2.6225 ;
      RECT  6.525 2.6225 18.2 5.0925 ;
      RECT  0.14 5.0925 5.825 7.085 ;
      RECT  6.525 5.0925 18.2 7.085 ;
      RECT  1.1075 7.085 5.825 12.47 ;
      RECT  6.525 7.085 18.2 12.47 ;
      RECT  6.525 12.47 18.2 17.665 ;
      RECT  5.825 18.1425 6.525 20.6125 ;
      RECT  6.525 17.665 18.2 18.1425 ;
      RECT  6.525 18.1425 18.2 20.6125 ;
      RECT  1.1075 20.6125 2.47 23.2925 ;
      RECT  3.17 20.6125 18.2 23.2925 ;
      RECT  1.1075 35.4325 2.47 35.465 ;
      RECT  1.1075 35.465 2.47 47.2125 ;
      RECT  2.47 35.465 3.17 47.2125 ;
      RECT  3.17 35.4325 15.48 35.465 ;
      RECT  3.17 35.465 15.48 47.2125 ;
      RECT  1.1075 23.2925 2.47 35.4325 ;
      RECT  3.17 23.2925 25.2 35.4325 ;
      RECT  1.1075 12.47 2.47 12.5025 ;
      RECT  1.1075 12.5025 2.47 17.665 ;
      RECT  2.47 12.47 3.17 12.5025 ;
      RECT  3.17 12.47 5.825 12.5025 ;
      RECT  3.17 12.5025 5.825 17.665 ;
      RECT  1.1075 17.665 2.47 18.1425 ;
      RECT  3.17 17.665 5.825 18.1425 ;
      RECT  1.1075 18.1425 2.47 20.6125 ;
      RECT  3.17 18.1425 5.825 20.6125 ;
   END
END    Ram_256_words
END    LIBRARY
